
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h1aa0d992;
    ram_cell[       1] = 32'h0;  // 32'h890cd40a;
    ram_cell[       2] = 32'h0;  // 32'h51ed81a5;
    ram_cell[       3] = 32'h0;  // 32'h7ced3dca;
    ram_cell[       4] = 32'h0;  // 32'hb2d586fd;
    ram_cell[       5] = 32'h0;  // 32'h5fa726fe;
    ram_cell[       6] = 32'h0;  // 32'h51c83745;
    ram_cell[       7] = 32'h0;  // 32'ha2664f45;
    ram_cell[       8] = 32'h0;  // 32'h72f962ab;
    ram_cell[       9] = 32'h0;  // 32'h8f90e5b9;
    ram_cell[      10] = 32'h0;  // 32'h1fa9177f;
    ram_cell[      11] = 32'h0;  // 32'hc5181ccd;
    ram_cell[      12] = 32'h0;  // 32'hfd6e73ec;
    ram_cell[      13] = 32'h0;  // 32'h37800ad8;
    ram_cell[      14] = 32'h0;  // 32'h0e918535;
    ram_cell[      15] = 32'h0;  // 32'h598af9d0;
    ram_cell[      16] = 32'h0;  // 32'h119efb03;
    ram_cell[      17] = 32'h0;  // 32'h54bd2cbc;
    ram_cell[      18] = 32'h0;  // 32'hc9bb7cca;
    ram_cell[      19] = 32'h0;  // 32'h5fbfc44a;
    ram_cell[      20] = 32'h0;  // 32'haf6744a4;
    ram_cell[      21] = 32'h0;  // 32'h971e7ca0;
    ram_cell[      22] = 32'h0;  // 32'h76eec5f4;
    ram_cell[      23] = 32'h0;  // 32'h5b3fd5d8;
    ram_cell[      24] = 32'h0;  // 32'hd2f0d355;
    ram_cell[      25] = 32'h0;  // 32'h6e04ad19;
    ram_cell[      26] = 32'h0;  // 32'ha8b83f0e;
    ram_cell[      27] = 32'h0;  // 32'hc97417c5;
    ram_cell[      28] = 32'h0;  // 32'hd7dbe210;
    ram_cell[      29] = 32'h0;  // 32'h72275a87;
    ram_cell[      30] = 32'h0;  // 32'h11b0ed60;
    ram_cell[      31] = 32'h0;  // 32'h5f26ba81;
    ram_cell[      32] = 32'h0;  // 32'h9610e1e6;
    ram_cell[      33] = 32'h0;  // 32'h26b0d849;
    ram_cell[      34] = 32'h0;  // 32'h39f76bb7;
    ram_cell[      35] = 32'h0;  // 32'h3614b31e;
    ram_cell[      36] = 32'h0;  // 32'h70945a9c;
    ram_cell[      37] = 32'h0;  // 32'he8bd6477;
    ram_cell[      38] = 32'h0;  // 32'h682884aa;
    ram_cell[      39] = 32'h0;  // 32'h371c149f;
    ram_cell[      40] = 32'h0;  // 32'hfe4286c7;
    ram_cell[      41] = 32'h0;  // 32'h8e99ab26;
    ram_cell[      42] = 32'h0;  // 32'h81109197;
    ram_cell[      43] = 32'h0;  // 32'h9b51266e;
    ram_cell[      44] = 32'h0;  // 32'h87ad03b8;
    ram_cell[      45] = 32'h0;  // 32'h9af67fe3;
    ram_cell[      46] = 32'h0;  // 32'h8607deaa;
    ram_cell[      47] = 32'h0;  // 32'h104a28c1;
    ram_cell[      48] = 32'h0;  // 32'h44c0835d;
    ram_cell[      49] = 32'h0;  // 32'h27db07f1;
    ram_cell[      50] = 32'h0;  // 32'h89581ff0;
    ram_cell[      51] = 32'h0;  // 32'ha4503784;
    ram_cell[      52] = 32'h0;  // 32'hbf4e21e3;
    ram_cell[      53] = 32'h0;  // 32'h45fd3abc;
    ram_cell[      54] = 32'h0;  // 32'hf95f6f29;
    ram_cell[      55] = 32'h0;  // 32'h6d337972;
    ram_cell[      56] = 32'h0;  // 32'he9cb1883;
    ram_cell[      57] = 32'h0;  // 32'hf50c1f45;
    ram_cell[      58] = 32'h0;  // 32'h973a8ea6;
    ram_cell[      59] = 32'h0;  // 32'h3b3c4838;
    ram_cell[      60] = 32'h0;  // 32'h48f1b5ef;
    ram_cell[      61] = 32'h0;  // 32'h6e3dfac9;
    ram_cell[      62] = 32'h0;  // 32'h95734a69;
    ram_cell[      63] = 32'h0;  // 32'h60a458b9;
    ram_cell[      64] = 32'h0;  // 32'h75951064;
    ram_cell[      65] = 32'h0;  // 32'h831313e2;
    ram_cell[      66] = 32'h0;  // 32'h9c19da55;
    ram_cell[      67] = 32'h0;  // 32'h181e3e19;
    ram_cell[      68] = 32'h0;  // 32'h8d0cdb77;
    ram_cell[      69] = 32'h0;  // 32'h1719f1a7;
    ram_cell[      70] = 32'h0;  // 32'h5a1eb6f3;
    ram_cell[      71] = 32'h0;  // 32'h4b2a1098;
    ram_cell[      72] = 32'h0;  // 32'he9651698;
    ram_cell[      73] = 32'h0;  // 32'hb8c291f5;
    ram_cell[      74] = 32'h0;  // 32'h41f804a3;
    ram_cell[      75] = 32'h0;  // 32'h012817c0;
    ram_cell[      76] = 32'h0;  // 32'h176eafdd;
    ram_cell[      77] = 32'h0;  // 32'hec614ca7;
    ram_cell[      78] = 32'h0;  // 32'hab99d821;
    ram_cell[      79] = 32'h0;  // 32'hac5a1f36;
    ram_cell[      80] = 32'h0;  // 32'h6ca96547;
    ram_cell[      81] = 32'h0;  // 32'hc083ff73;
    ram_cell[      82] = 32'h0;  // 32'h2356ea4b;
    ram_cell[      83] = 32'h0;  // 32'h93034896;
    ram_cell[      84] = 32'h0;  // 32'hf9765ba2;
    ram_cell[      85] = 32'h0;  // 32'h90f3cb11;
    ram_cell[      86] = 32'h0;  // 32'h2ea06600;
    ram_cell[      87] = 32'h0;  // 32'h9d5f5d62;
    ram_cell[      88] = 32'h0;  // 32'h1fea052b;
    ram_cell[      89] = 32'h0;  // 32'h7b82b3e1;
    ram_cell[      90] = 32'h0;  // 32'h1d6de7a3;
    ram_cell[      91] = 32'h0;  // 32'h0446b861;
    ram_cell[      92] = 32'h0;  // 32'h37d25453;
    ram_cell[      93] = 32'h0;  // 32'h28b34d4d;
    ram_cell[      94] = 32'h0;  // 32'h924084cb;
    ram_cell[      95] = 32'h0;  // 32'hb5ab8513;
    ram_cell[      96] = 32'h0;  // 32'h95414d7f;
    ram_cell[      97] = 32'h0;  // 32'hfa343cf4;
    ram_cell[      98] = 32'h0;  // 32'hd5b9dcd2;
    ram_cell[      99] = 32'h0;  // 32'h31ab12fd;
    ram_cell[     100] = 32'h0;  // 32'h1a3fa41c;
    ram_cell[     101] = 32'h0;  // 32'h702996d6;
    ram_cell[     102] = 32'h0;  // 32'h4967817e;
    ram_cell[     103] = 32'h0;  // 32'hcfd12cdf;
    ram_cell[     104] = 32'h0;  // 32'ha1789d35;
    ram_cell[     105] = 32'h0;  // 32'hf370a4cf;
    ram_cell[     106] = 32'h0;  // 32'hce4bfd0a;
    ram_cell[     107] = 32'h0;  // 32'hdb8dfee7;
    ram_cell[     108] = 32'h0;  // 32'hb594212c;
    ram_cell[     109] = 32'h0;  // 32'h7b4089e2;
    ram_cell[     110] = 32'h0;  // 32'h14115c7f;
    ram_cell[     111] = 32'h0;  // 32'h69595296;
    ram_cell[     112] = 32'h0;  // 32'haf1a5211;
    ram_cell[     113] = 32'h0;  // 32'hcd4f80bf;
    ram_cell[     114] = 32'h0;  // 32'hb982edf7;
    ram_cell[     115] = 32'h0;  // 32'h1d0230c8;
    ram_cell[     116] = 32'h0;  // 32'h05de391c;
    ram_cell[     117] = 32'h0;  // 32'h824dee21;
    ram_cell[     118] = 32'h0;  // 32'h98fe79aa;
    ram_cell[     119] = 32'h0;  // 32'h7569dfb7;
    ram_cell[     120] = 32'h0;  // 32'hf30df688;
    ram_cell[     121] = 32'h0;  // 32'hf197a90a;
    ram_cell[     122] = 32'h0;  // 32'h3a4757c1;
    ram_cell[     123] = 32'h0;  // 32'h1984486e;
    ram_cell[     124] = 32'h0;  // 32'h108bcf94;
    ram_cell[     125] = 32'h0;  // 32'hcca634fb;
    ram_cell[     126] = 32'h0;  // 32'h9e8e7483;
    ram_cell[     127] = 32'h0;  // 32'hd4d2dd60;
    ram_cell[     128] = 32'h0;  // 32'he31305c1;
    ram_cell[     129] = 32'h0;  // 32'h31b28e43;
    ram_cell[     130] = 32'h0;  // 32'h6b242501;
    ram_cell[     131] = 32'h0;  // 32'h7cf21f4f;
    ram_cell[     132] = 32'h0;  // 32'hcfac26d2;
    ram_cell[     133] = 32'h0;  // 32'h9eef6f32;
    ram_cell[     134] = 32'h0;  // 32'haebdca0d;
    ram_cell[     135] = 32'h0;  // 32'hd24f5551;
    ram_cell[     136] = 32'h0;  // 32'hc29cf3f6;
    ram_cell[     137] = 32'h0;  // 32'ha2d4b01f;
    ram_cell[     138] = 32'h0;  // 32'hfbb9c3f1;
    ram_cell[     139] = 32'h0;  // 32'h161ee364;
    ram_cell[     140] = 32'h0;  // 32'h72ca6eb5;
    ram_cell[     141] = 32'h0;  // 32'h444c6445;
    ram_cell[     142] = 32'h0;  // 32'haabe744a;
    ram_cell[     143] = 32'h0;  // 32'h25367ec2;
    ram_cell[     144] = 32'h0;  // 32'h03a96f1a;
    ram_cell[     145] = 32'h0;  // 32'hd36a2b77;
    ram_cell[     146] = 32'h0;  // 32'hf9e164e8;
    ram_cell[     147] = 32'h0;  // 32'h5996ac1c;
    ram_cell[     148] = 32'h0;  // 32'h794b1ef7;
    ram_cell[     149] = 32'h0;  // 32'hd23cdf90;
    ram_cell[     150] = 32'h0;  // 32'hdc938c37;
    ram_cell[     151] = 32'h0;  // 32'h7e0f5af6;
    ram_cell[     152] = 32'h0;  // 32'hc32bdc8d;
    ram_cell[     153] = 32'h0;  // 32'hf71798c4;
    ram_cell[     154] = 32'h0;  // 32'he3f4b0e1;
    ram_cell[     155] = 32'h0;  // 32'h313c27a4;
    ram_cell[     156] = 32'h0;  // 32'h736dbf22;
    ram_cell[     157] = 32'h0;  // 32'h1f7676fa;
    ram_cell[     158] = 32'h0;  // 32'h3c26d9a8;
    ram_cell[     159] = 32'h0;  // 32'he36bb9bf;
    ram_cell[     160] = 32'h0;  // 32'h9bd8c7d3;
    ram_cell[     161] = 32'h0;  // 32'ha28ec1be;
    ram_cell[     162] = 32'h0;  // 32'h5996a382;
    ram_cell[     163] = 32'h0;  // 32'h3188bca0;
    ram_cell[     164] = 32'h0;  // 32'hc1d415ea;
    ram_cell[     165] = 32'h0;  // 32'hb8e3683c;
    ram_cell[     166] = 32'h0;  // 32'h4c95200b;
    ram_cell[     167] = 32'h0;  // 32'hcb6de470;
    ram_cell[     168] = 32'h0;  // 32'h212fe2ca;
    ram_cell[     169] = 32'h0;  // 32'hd56cb46b;
    ram_cell[     170] = 32'h0;  // 32'h87df24a7;
    ram_cell[     171] = 32'h0;  // 32'h5ead63ee;
    ram_cell[     172] = 32'h0;  // 32'h3dfefafc;
    ram_cell[     173] = 32'h0;  // 32'h18335dec;
    ram_cell[     174] = 32'h0;  // 32'h61631dc9;
    ram_cell[     175] = 32'h0;  // 32'hecc7e28e;
    ram_cell[     176] = 32'h0;  // 32'h20cb1273;
    ram_cell[     177] = 32'h0;  // 32'h817628f1;
    ram_cell[     178] = 32'h0;  // 32'h36db43e6;
    ram_cell[     179] = 32'h0;  // 32'h4f32003a;
    ram_cell[     180] = 32'h0;  // 32'hf83a34ca;
    ram_cell[     181] = 32'h0;  // 32'h873b55d9;
    ram_cell[     182] = 32'h0;  // 32'he67b1f60;
    ram_cell[     183] = 32'h0;  // 32'h533a4d6a;
    ram_cell[     184] = 32'h0;  // 32'h139b55db;
    ram_cell[     185] = 32'h0;  // 32'hfa20fa57;
    ram_cell[     186] = 32'h0;  // 32'h13905bd8;
    ram_cell[     187] = 32'h0;  // 32'h9a880ba0;
    ram_cell[     188] = 32'h0;  // 32'h8a801421;
    ram_cell[     189] = 32'h0;  // 32'hf923bbbe;
    ram_cell[     190] = 32'h0;  // 32'h3662d354;
    ram_cell[     191] = 32'h0;  // 32'h95327942;
    ram_cell[     192] = 32'h0;  // 32'h683d110a;
    ram_cell[     193] = 32'h0;  // 32'haef0c7fe;
    ram_cell[     194] = 32'h0;  // 32'h04509260;
    ram_cell[     195] = 32'h0;  // 32'h363b10d1;
    ram_cell[     196] = 32'h0;  // 32'hd1ba7915;
    ram_cell[     197] = 32'h0;  // 32'hf034dc40;
    ram_cell[     198] = 32'h0;  // 32'h94408e01;
    ram_cell[     199] = 32'h0;  // 32'hc25a9f29;
    ram_cell[     200] = 32'h0;  // 32'ha30bf09b;
    ram_cell[     201] = 32'h0;  // 32'h6582b120;
    ram_cell[     202] = 32'h0;  // 32'h798e40db;
    ram_cell[     203] = 32'h0;  // 32'h9c331aa1;
    ram_cell[     204] = 32'h0;  // 32'hbf80c37d;
    ram_cell[     205] = 32'h0;  // 32'hfd120866;
    ram_cell[     206] = 32'h0;  // 32'h233d8638;
    ram_cell[     207] = 32'h0;  // 32'h3e300e1b;
    ram_cell[     208] = 32'h0;  // 32'h58303843;
    ram_cell[     209] = 32'h0;  // 32'he9a04d94;
    ram_cell[     210] = 32'h0;  // 32'hdf5019ec;
    ram_cell[     211] = 32'h0;  // 32'h2b300dfa;
    ram_cell[     212] = 32'h0;  // 32'ha255477e;
    ram_cell[     213] = 32'h0;  // 32'h9a21d51e;
    ram_cell[     214] = 32'h0;  // 32'h0b5e7514;
    ram_cell[     215] = 32'h0;  // 32'h1b0c0bb7;
    ram_cell[     216] = 32'h0;  // 32'hac0c06a6;
    ram_cell[     217] = 32'h0;  // 32'h1cde7def;
    ram_cell[     218] = 32'h0;  // 32'h8c8133ab;
    ram_cell[     219] = 32'h0;  // 32'h2fb3227d;
    ram_cell[     220] = 32'h0;  // 32'hffef8d08;
    ram_cell[     221] = 32'h0;  // 32'h30573f12;
    ram_cell[     222] = 32'h0;  // 32'h37070494;
    ram_cell[     223] = 32'h0;  // 32'h46284415;
    ram_cell[     224] = 32'h0;  // 32'hb7d39d45;
    ram_cell[     225] = 32'h0;  // 32'h5434c783;
    ram_cell[     226] = 32'h0;  // 32'hbf213faa;
    ram_cell[     227] = 32'h0;  // 32'h1637b851;
    ram_cell[     228] = 32'h0;  // 32'ha453d5a2;
    ram_cell[     229] = 32'h0;  // 32'h94de7c10;
    ram_cell[     230] = 32'h0;  // 32'h8ed7beb1;
    ram_cell[     231] = 32'h0;  // 32'hcf13a08b;
    ram_cell[     232] = 32'h0;  // 32'h61aeb632;
    ram_cell[     233] = 32'h0;  // 32'h69dee95c;
    ram_cell[     234] = 32'h0;  // 32'he3e39f37;
    ram_cell[     235] = 32'h0;  // 32'hdb614fde;
    ram_cell[     236] = 32'h0;  // 32'hb20b1624;
    ram_cell[     237] = 32'h0;  // 32'h264fc98d;
    ram_cell[     238] = 32'h0;  // 32'h41af245d;
    ram_cell[     239] = 32'h0;  // 32'h1ebcafa4;
    ram_cell[     240] = 32'h0;  // 32'he24e2660;
    ram_cell[     241] = 32'h0;  // 32'hc6c19588;
    ram_cell[     242] = 32'h0;  // 32'h66a011a0;
    ram_cell[     243] = 32'h0;  // 32'he049f103;
    ram_cell[     244] = 32'h0;  // 32'hd58e742d;
    ram_cell[     245] = 32'h0;  // 32'h263fbf1f;
    ram_cell[     246] = 32'h0;  // 32'hac3efbf0;
    ram_cell[     247] = 32'h0;  // 32'h3f6951a4;
    ram_cell[     248] = 32'h0;  // 32'hf7c4d297;
    ram_cell[     249] = 32'h0;  // 32'h1acb5d91;
    ram_cell[     250] = 32'h0;  // 32'h91c4a437;
    ram_cell[     251] = 32'h0;  // 32'h114ecc44;
    ram_cell[     252] = 32'h0;  // 32'hc79f915b;
    ram_cell[     253] = 32'h0;  // 32'hbe557ef6;
    ram_cell[     254] = 32'h0;  // 32'hb494a1e9;
    ram_cell[     255] = 32'h0;  // 32'h178b0418;
    // src matrix A
    ram_cell[     256] = 32'h0574d8e9;
    ram_cell[     257] = 32'h7995cb8e;
    ram_cell[     258] = 32'hf64f3b79;
    ram_cell[     259] = 32'h55cb7f87;
    ram_cell[     260] = 32'hd89ac3c5;
    ram_cell[     261] = 32'h5bca3c15;
    ram_cell[     262] = 32'h237dfe40;
    ram_cell[     263] = 32'hb8845115;
    ram_cell[     264] = 32'hb32426e6;
    ram_cell[     265] = 32'h9badd8d7;
    ram_cell[     266] = 32'h0ceb9ece;
    ram_cell[     267] = 32'h0ca459f4;
    ram_cell[     268] = 32'h869924f4;
    ram_cell[     269] = 32'h8e8d0db3;
    ram_cell[     270] = 32'h1fb24328;
    ram_cell[     271] = 32'haa328cec;
    ram_cell[     272] = 32'hc7c1a770;
    ram_cell[     273] = 32'ha9f66859;
    ram_cell[     274] = 32'hce2a91f8;
    ram_cell[     275] = 32'hbe3d31e6;
    ram_cell[     276] = 32'h77708f74;
    ram_cell[     277] = 32'h7531ec5d;
    ram_cell[     278] = 32'h9cf35df4;
    ram_cell[     279] = 32'h7326987c;
    ram_cell[     280] = 32'h159f5224;
    ram_cell[     281] = 32'h4175f110;
    ram_cell[     282] = 32'ha549888f;
    ram_cell[     283] = 32'he83a78c3;
    ram_cell[     284] = 32'hb0598797;
    ram_cell[     285] = 32'hd26fe7e1;
    ram_cell[     286] = 32'h624840aa;
    ram_cell[     287] = 32'h7f86b50e;
    ram_cell[     288] = 32'hfb861e2e;
    ram_cell[     289] = 32'haad401bd;
    ram_cell[     290] = 32'hd1b49ea8;
    ram_cell[     291] = 32'ha3ca9839;
    ram_cell[     292] = 32'he47982fe;
    ram_cell[     293] = 32'h7ad0659c;
    ram_cell[     294] = 32'h27ed4702;
    ram_cell[     295] = 32'h6410d655;
    ram_cell[     296] = 32'h780ef93e;
    ram_cell[     297] = 32'hbac9ca4d;
    ram_cell[     298] = 32'h41531f04;
    ram_cell[     299] = 32'h9fe81d2e;
    ram_cell[     300] = 32'hbf8c919f;
    ram_cell[     301] = 32'h17a21ddf;
    ram_cell[     302] = 32'h7ba6bb3c;
    ram_cell[     303] = 32'h047495d5;
    ram_cell[     304] = 32'h5923a8a0;
    ram_cell[     305] = 32'he38f3e42;
    ram_cell[     306] = 32'ha8b7f468;
    ram_cell[     307] = 32'hc66756a6;
    ram_cell[     308] = 32'h9e71fc2a;
    ram_cell[     309] = 32'h73e6901f;
    ram_cell[     310] = 32'h49f6dd15;
    ram_cell[     311] = 32'he576ac43;
    ram_cell[     312] = 32'h78311e53;
    ram_cell[     313] = 32'h9d15592e;
    ram_cell[     314] = 32'h31540d29;
    ram_cell[     315] = 32'hc45cdb10;
    ram_cell[     316] = 32'h2f2558c5;
    ram_cell[     317] = 32'hb282a3ef;
    ram_cell[     318] = 32'h79e207db;
    ram_cell[     319] = 32'he3986802;
    ram_cell[     320] = 32'hb175f1ab;
    ram_cell[     321] = 32'h0d32a5ef;
    ram_cell[     322] = 32'hdad68c38;
    ram_cell[     323] = 32'hec1131c9;
    ram_cell[     324] = 32'h2121d832;
    ram_cell[     325] = 32'h69909796;
    ram_cell[     326] = 32'h8f8554a7;
    ram_cell[     327] = 32'h77be00a3;
    ram_cell[     328] = 32'h904abceb;
    ram_cell[     329] = 32'h69d2adf5;
    ram_cell[     330] = 32'hf30d67f2;
    ram_cell[     331] = 32'h0cba0435;
    ram_cell[     332] = 32'h7f5ab317;
    ram_cell[     333] = 32'h4bb04db3;
    ram_cell[     334] = 32'h52b9b84b;
    ram_cell[     335] = 32'he60946c6;
    ram_cell[     336] = 32'hde5daafa;
    ram_cell[     337] = 32'h0d02354d;
    ram_cell[     338] = 32'h83acd3e2;
    ram_cell[     339] = 32'h52fb47fb;
    ram_cell[     340] = 32'hcd9a6e06;
    ram_cell[     341] = 32'ha6fc8237;
    ram_cell[     342] = 32'hdb6ea682;
    ram_cell[     343] = 32'hc2ed2de8;
    ram_cell[     344] = 32'he60aa70d;
    ram_cell[     345] = 32'h0b953cb8;
    ram_cell[     346] = 32'h15575969;
    ram_cell[     347] = 32'h1318b60a;
    ram_cell[     348] = 32'hd902fa78;
    ram_cell[     349] = 32'hc74fb734;
    ram_cell[     350] = 32'h081b2b57;
    ram_cell[     351] = 32'ha79a9e13;
    ram_cell[     352] = 32'h222a22eb;
    ram_cell[     353] = 32'hfd3b87de;
    ram_cell[     354] = 32'ha93735f3;
    ram_cell[     355] = 32'h6737effa;
    ram_cell[     356] = 32'h01140585;
    ram_cell[     357] = 32'h0500002d;
    ram_cell[     358] = 32'h3e43aeb4;
    ram_cell[     359] = 32'h4587117f;
    ram_cell[     360] = 32'h963e526d;
    ram_cell[     361] = 32'hd1f853a9;
    ram_cell[     362] = 32'hadd78021;
    ram_cell[     363] = 32'h3ddaa5df;
    ram_cell[     364] = 32'h82fb762e;
    ram_cell[     365] = 32'h6b687c27;
    ram_cell[     366] = 32'hd3284bfe;
    ram_cell[     367] = 32'hb2c4a55f;
    ram_cell[     368] = 32'h9b664c1b;
    ram_cell[     369] = 32'h05c9c7d4;
    ram_cell[     370] = 32'h0f99db03;
    ram_cell[     371] = 32'h17f81df5;
    ram_cell[     372] = 32'hc2d198bf;
    ram_cell[     373] = 32'h130d9b5e;
    ram_cell[     374] = 32'h87cd0948;
    ram_cell[     375] = 32'haf4e033b;
    ram_cell[     376] = 32'h2acc34bd;
    ram_cell[     377] = 32'hbd6377d2;
    ram_cell[     378] = 32'hd69cbb66;
    ram_cell[     379] = 32'h2644780f;
    ram_cell[     380] = 32'h488d1bbe;
    ram_cell[     381] = 32'h0fd23f3f;
    ram_cell[     382] = 32'h06fbb913;
    ram_cell[     383] = 32'h3474c537;
    ram_cell[     384] = 32'hfdb4d384;
    ram_cell[     385] = 32'h8e4550fd;
    ram_cell[     386] = 32'h4cac543a;
    ram_cell[     387] = 32'h1b8cf89d;
    ram_cell[     388] = 32'h173d7fdf;
    ram_cell[     389] = 32'h4ffbec67;
    ram_cell[     390] = 32'hef1b471c;
    ram_cell[     391] = 32'hda3fd801;
    ram_cell[     392] = 32'h1bd0112f;
    ram_cell[     393] = 32'h93e461da;
    ram_cell[     394] = 32'h2d5fc1ed;
    ram_cell[     395] = 32'h9f6ca179;
    ram_cell[     396] = 32'h3b08330d;
    ram_cell[     397] = 32'h0f8fdaf0;
    ram_cell[     398] = 32'h038aa522;
    ram_cell[     399] = 32'h79008019;
    ram_cell[     400] = 32'h3ded5927;
    ram_cell[     401] = 32'hd6477bc1;
    ram_cell[     402] = 32'he5c03ade;
    ram_cell[     403] = 32'ha954f5d6;
    ram_cell[     404] = 32'hdf6777dc;
    ram_cell[     405] = 32'h7f58d482;
    ram_cell[     406] = 32'hcfa43fe3;
    ram_cell[     407] = 32'h964322fd;
    ram_cell[     408] = 32'h9780fb9e;
    ram_cell[     409] = 32'hfdd350b3;
    ram_cell[     410] = 32'h7b089a1d;
    ram_cell[     411] = 32'hdc311a55;
    ram_cell[     412] = 32'h80b05258;
    ram_cell[     413] = 32'h258a1f9a;
    ram_cell[     414] = 32'h39f2bfc7;
    ram_cell[     415] = 32'h23af139f;
    ram_cell[     416] = 32'h628751c7;
    ram_cell[     417] = 32'h111fdd8e;
    ram_cell[     418] = 32'ha1374d2b;
    ram_cell[     419] = 32'h90bd04c3;
    ram_cell[     420] = 32'h59fc75ec;
    ram_cell[     421] = 32'h600b6f2d;
    ram_cell[     422] = 32'h1aefbb0e;
    ram_cell[     423] = 32'hc0553c2b;
    ram_cell[     424] = 32'h7f292d95;
    ram_cell[     425] = 32'h00f7608f;
    ram_cell[     426] = 32'h6ce4eff2;
    ram_cell[     427] = 32'h9dba84ad;
    ram_cell[     428] = 32'h199aa5b2;
    ram_cell[     429] = 32'h3650531f;
    ram_cell[     430] = 32'he40f442d;
    ram_cell[     431] = 32'h11fd2ec8;
    ram_cell[     432] = 32'h69394b5b;
    ram_cell[     433] = 32'h39a73fc0;
    ram_cell[     434] = 32'h01dfd546;
    ram_cell[     435] = 32'h2eeb5cd7;
    ram_cell[     436] = 32'hde68257b;
    ram_cell[     437] = 32'hccf5a0f2;
    ram_cell[     438] = 32'h5a76edaa;
    ram_cell[     439] = 32'h54e4ab29;
    ram_cell[     440] = 32'h750618e3;
    ram_cell[     441] = 32'h81661fa6;
    ram_cell[     442] = 32'he2a3e416;
    ram_cell[     443] = 32'hb219d125;
    ram_cell[     444] = 32'ha30edd1a;
    ram_cell[     445] = 32'he0e79833;
    ram_cell[     446] = 32'hba1e7d9f;
    ram_cell[     447] = 32'h55f4d990;
    ram_cell[     448] = 32'h00cbff78;
    ram_cell[     449] = 32'h57f694a6;
    ram_cell[     450] = 32'hefceb2f2;
    ram_cell[     451] = 32'he1d7209b;
    ram_cell[     452] = 32'h02c1acef;
    ram_cell[     453] = 32'ha7f5c73b;
    ram_cell[     454] = 32'hd89f7865;
    ram_cell[     455] = 32'hcf5582b9;
    ram_cell[     456] = 32'h9576a27a;
    ram_cell[     457] = 32'h4a6cdd92;
    ram_cell[     458] = 32'haac5b23b;
    ram_cell[     459] = 32'h1a133719;
    ram_cell[     460] = 32'h60dd93e2;
    ram_cell[     461] = 32'hc9f6386d;
    ram_cell[     462] = 32'h88aceffe;
    ram_cell[     463] = 32'h8d7c9fb0;
    ram_cell[     464] = 32'h94739e70;
    ram_cell[     465] = 32'h2ec659c6;
    ram_cell[     466] = 32'h2ebea950;
    ram_cell[     467] = 32'h14331bae;
    ram_cell[     468] = 32'h448294ca;
    ram_cell[     469] = 32'h68da3ac3;
    ram_cell[     470] = 32'h39a96da5;
    ram_cell[     471] = 32'hf2a8f2b8;
    ram_cell[     472] = 32'hed58f02e;
    ram_cell[     473] = 32'hf28d3382;
    ram_cell[     474] = 32'h123b14f7;
    ram_cell[     475] = 32'h9727019e;
    ram_cell[     476] = 32'h5c37916f;
    ram_cell[     477] = 32'h6f6ead51;
    ram_cell[     478] = 32'h746b58d7;
    ram_cell[     479] = 32'h387b7f0b;
    ram_cell[     480] = 32'h59a7b85c;
    ram_cell[     481] = 32'h5a623182;
    ram_cell[     482] = 32'hbb7cd341;
    ram_cell[     483] = 32'hc582009f;
    ram_cell[     484] = 32'h88d9c139;
    ram_cell[     485] = 32'h041db4ff;
    ram_cell[     486] = 32'hdbd42a99;
    ram_cell[     487] = 32'h1867b9b5;
    ram_cell[     488] = 32'h05333483;
    ram_cell[     489] = 32'h439c3832;
    ram_cell[     490] = 32'h7ce2c80b;
    ram_cell[     491] = 32'hfe43d99c;
    ram_cell[     492] = 32'h4e70573f;
    ram_cell[     493] = 32'h0983c962;
    ram_cell[     494] = 32'h6a03666d;
    ram_cell[     495] = 32'hfe5510c3;
    ram_cell[     496] = 32'hc9b60b50;
    ram_cell[     497] = 32'h3883acbb;
    ram_cell[     498] = 32'h556efe80;
    ram_cell[     499] = 32'h017bb76a;
    ram_cell[     500] = 32'h9a46f9f2;
    ram_cell[     501] = 32'hf5043486;
    ram_cell[     502] = 32'h81a33ba1;
    ram_cell[     503] = 32'h7200782c;
    ram_cell[     504] = 32'h2d556c54;
    ram_cell[     505] = 32'hcdd40e7a;
    ram_cell[     506] = 32'h5ee5ce62;
    ram_cell[     507] = 32'hb1fd61d1;
    ram_cell[     508] = 32'hf2a87e07;
    ram_cell[     509] = 32'h515f33a1;
    ram_cell[     510] = 32'h7f89d1a7;
    ram_cell[     511] = 32'hafb13dea;
    // src matrix B
    ram_cell[     512] = 32'hc11a5191;
    ram_cell[     513] = 32'hb9589512;
    ram_cell[     514] = 32'h78935c42;
    ram_cell[     515] = 32'hf86a452a;
    ram_cell[     516] = 32'h0655b141;
    ram_cell[     517] = 32'hd258caf8;
    ram_cell[     518] = 32'hf3eb86fc;
    ram_cell[     519] = 32'h1f7f46e8;
    ram_cell[     520] = 32'h244cb162;
    ram_cell[     521] = 32'ha2a85df5;
    ram_cell[     522] = 32'h70d399ca;
    ram_cell[     523] = 32'h20b19e7c;
    ram_cell[     524] = 32'h5748dd87;
    ram_cell[     525] = 32'h424d7278;
    ram_cell[     526] = 32'h6e8553c2;
    ram_cell[     527] = 32'h63fe9733;
    ram_cell[     528] = 32'h55f265ea;
    ram_cell[     529] = 32'h0a1d87c4;
    ram_cell[     530] = 32'h15723316;
    ram_cell[     531] = 32'ha0f6bccd;
    ram_cell[     532] = 32'h303ba057;
    ram_cell[     533] = 32'hd1f8fb64;
    ram_cell[     534] = 32'h2cfebf7a;
    ram_cell[     535] = 32'h6fb4723f;
    ram_cell[     536] = 32'h47ded4aa;
    ram_cell[     537] = 32'hca2a484a;
    ram_cell[     538] = 32'hc440582b;
    ram_cell[     539] = 32'hf02e682e;
    ram_cell[     540] = 32'hf18db90c;
    ram_cell[     541] = 32'h0198378a;
    ram_cell[     542] = 32'hf2d5d63a;
    ram_cell[     543] = 32'h1dba0879;
    ram_cell[     544] = 32'hbbcf2d00;
    ram_cell[     545] = 32'h27c7e1f8;
    ram_cell[     546] = 32'h82334af0;
    ram_cell[     547] = 32'h3c75afae;
    ram_cell[     548] = 32'h37fcd593;
    ram_cell[     549] = 32'h0d358e89;
    ram_cell[     550] = 32'h9af43e51;
    ram_cell[     551] = 32'ha37dbd9f;
    ram_cell[     552] = 32'hf259108b;
    ram_cell[     553] = 32'hb83ace95;
    ram_cell[     554] = 32'hcef4305d;
    ram_cell[     555] = 32'hd824e160;
    ram_cell[     556] = 32'h0dc94f23;
    ram_cell[     557] = 32'ha88777f6;
    ram_cell[     558] = 32'h0aa66d1b;
    ram_cell[     559] = 32'h8f0dd393;
    ram_cell[     560] = 32'h32a104d3;
    ram_cell[     561] = 32'ha730a9fe;
    ram_cell[     562] = 32'hf311b5e7;
    ram_cell[     563] = 32'hc6351a2e;
    ram_cell[     564] = 32'h90f0de56;
    ram_cell[     565] = 32'h141a722c;
    ram_cell[     566] = 32'h9c8ada5f;
    ram_cell[     567] = 32'hc454edff;
    ram_cell[     568] = 32'hb061f6a4;
    ram_cell[     569] = 32'ha1498d73;
    ram_cell[     570] = 32'hf6caf6ba;
    ram_cell[     571] = 32'h6ca534f9;
    ram_cell[     572] = 32'h4ce6fac5;
    ram_cell[     573] = 32'h14245b7d;
    ram_cell[     574] = 32'h150445b3;
    ram_cell[     575] = 32'h0b78546a;
    ram_cell[     576] = 32'h1ceaceba;
    ram_cell[     577] = 32'h04cc5d23;
    ram_cell[     578] = 32'h0ba331d5;
    ram_cell[     579] = 32'h7e61b9cd;
    ram_cell[     580] = 32'h6163139c;
    ram_cell[     581] = 32'h3aaca620;
    ram_cell[     582] = 32'h07a4b427;
    ram_cell[     583] = 32'h2b87ab3d;
    ram_cell[     584] = 32'hea6f7b4b;
    ram_cell[     585] = 32'h97c1214c;
    ram_cell[     586] = 32'h31f72f43;
    ram_cell[     587] = 32'h206ea9aa;
    ram_cell[     588] = 32'h06a75489;
    ram_cell[     589] = 32'h23afe5c6;
    ram_cell[     590] = 32'h5cd1c2b9;
    ram_cell[     591] = 32'h6b600878;
    ram_cell[     592] = 32'he981251c;
    ram_cell[     593] = 32'h9a7cc5bf;
    ram_cell[     594] = 32'haf242f5e;
    ram_cell[     595] = 32'h2559d139;
    ram_cell[     596] = 32'hd6e346da;
    ram_cell[     597] = 32'h0bf94563;
    ram_cell[     598] = 32'hec87fec1;
    ram_cell[     599] = 32'h045a4a18;
    ram_cell[     600] = 32'hd0ac62bb;
    ram_cell[     601] = 32'h0a99adb1;
    ram_cell[     602] = 32'hd9de03f2;
    ram_cell[     603] = 32'hc27823c4;
    ram_cell[     604] = 32'h05bcafca;
    ram_cell[     605] = 32'ha0eb7a78;
    ram_cell[     606] = 32'hced797b7;
    ram_cell[     607] = 32'hec95094b;
    ram_cell[     608] = 32'h3ec28324;
    ram_cell[     609] = 32'h66014138;
    ram_cell[     610] = 32'he2874afb;
    ram_cell[     611] = 32'h11e902fc;
    ram_cell[     612] = 32'h0db9905c;
    ram_cell[     613] = 32'hd318a481;
    ram_cell[     614] = 32'hec16e887;
    ram_cell[     615] = 32'h77cc0257;
    ram_cell[     616] = 32'h8ad801b3;
    ram_cell[     617] = 32'h5cfe08c4;
    ram_cell[     618] = 32'he68066d1;
    ram_cell[     619] = 32'haf11c745;
    ram_cell[     620] = 32'h2caf40e1;
    ram_cell[     621] = 32'h8a4ccae9;
    ram_cell[     622] = 32'h3ae676ea;
    ram_cell[     623] = 32'h33e6821f;
    ram_cell[     624] = 32'he00bda1f;
    ram_cell[     625] = 32'h2ca43730;
    ram_cell[     626] = 32'h7aca26f9;
    ram_cell[     627] = 32'hdbd25204;
    ram_cell[     628] = 32'hfcb5707f;
    ram_cell[     629] = 32'he74aaa4f;
    ram_cell[     630] = 32'hb5008993;
    ram_cell[     631] = 32'h21ff5c4e;
    ram_cell[     632] = 32'h7bade74f;
    ram_cell[     633] = 32'h029073ce;
    ram_cell[     634] = 32'h8ec9c785;
    ram_cell[     635] = 32'h824f76fb;
    ram_cell[     636] = 32'h840f9b1f;
    ram_cell[     637] = 32'h5caaef57;
    ram_cell[     638] = 32'h18ec3c22;
    ram_cell[     639] = 32'h00143928;
    ram_cell[     640] = 32'hc0f0ec91;
    ram_cell[     641] = 32'ha449893f;
    ram_cell[     642] = 32'h9f7bebce;
    ram_cell[     643] = 32'he73d482c;
    ram_cell[     644] = 32'h1286d6e7;
    ram_cell[     645] = 32'hfa863b66;
    ram_cell[     646] = 32'h3e6aa80b;
    ram_cell[     647] = 32'h37f87969;
    ram_cell[     648] = 32'hee5e989e;
    ram_cell[     649] = 32'hd2bcb9fe;
    ram_cell[     650] = 32'h0fb14764;
    ram_cell[     651] = 32'h5c536250;
    ram_cell[     652] = 32'h2471daa2;
    ram_cell[     653] = 32'h8ffd0ab3;
    ram_cell[     654] = 32'hbaa9643d;
    ram_cell[     655] = 32'h16b036c3;
    ram_cell[     656] = 32'h2bbd8f64;
    ram_cell[     657] = 32'hfecda173;
    ram_cell[     658] = 32'h38a68e4f;
    ram_cell[     659] = 32'h034943a6;
    ram_cell[     660] = 32'h90f06d15;
    ram_cell[     661] = 32'hd5b66585;
    ram_cell[     662] = 32'he7742de4;
    ram_cell[     663] = 32'h03cc12a6;
    ram_cell[     664] = 32'h035aa93c;
    ram_cell[     665] = 32'hbf1c178e;
    ram_cell[     666] = 32'h06cc2475;
    ram_cell[     667] = 32'h12f43c6a;
    ram_cell[     668] = 32'hda0bbd6b;
    ram_cell[     669] = 32'h0e564890;
    ram_cell[     670] = 32'hef0fe040;
    ram_cell[     671] = 32'h17970932;
    ram_cell[     672] = 32'hb98e7392;
    ram_cell[     673] = 32'hef74eba8;
    ram_cell[     674] = 32'h29ac9e14;
    ram_cell[     675] = 32'h318c6b58;
    ram_cell[     676] = 32'h0d16155e;
    ram_cell[     677] = 32'h5ad3c036;
    ram_cell[     678] = 32'hcff4d676;
    ram_cell[     679] = 32'hec478967;
    ram_cell[     680] = 32'hf6ceb7bf;
    ram_cell[     681] = 32'heee11007;
    ram_cell[     682] = 32'h4c7efb84;
    ram_cell[     683] = 32'hbf5399d1;
    ram_cell[     684] = 32'h5d0a9055;
    ram_cell[     685] = 32'h9d1c4d40;
    ram_cell[     686] = 32'hfb9f534a;
    ram_cell[     687] = 32'h34e1363c;
    ram_cell[     688] = 32'h2368d381;
    ram_cell[     689] = 32'h6f073c9f;
    ram_cell[     690] = 32'h2edc3efb;
    ram_cell[     691] = 32'hf6618c69;
    ram_cell[     692] = 32'hb61c1615;
    ram_cell[     693] = 32'h5f35ba4d;
    ram_cell[     694] = 32'hcde1fdbc;
    ram_cell[     695] = 32'hd0f36231;
    ram_cell[     696] = 32'hcbc2fd01;
    ram_cell[     697] = 32'ha262cfae;
    ram_cell[     698] = 32'hf97f9f27;
    ram_cell[     699] = 32'h0b658374;
    ram_cell[     700] = 32'hddcf7af2;
    ram_cell[     701] = 32'h942e72a3;
    ram_cell[     702] = 32'h9d15e816;
    ram_cell[     703] = 32'hced842ba;
    ram_cell[     704] = 32'hc5389289;
    ram_cell[     705] = 32'h0b26aae7;
    ram_cell[     706] = 32'h46519ede;
    ram_cell[     707] = 32'h00e3b2a3;
    ram_cell[     708] = 32'h14abbaad;
    ram_cell[     709] = 32'h757fbb28;
    ram_cell[     710] = 32'hb1ad1ffd;
    ram_cell[     711] = 32'h3f83ddc1;
    ram_cell[     712] = 32'h5bda3a0d;
    ram_cell[     713] = 32'hb5f59e5e;
    ram_cell[     714] = 32'hced0a5ab;
    ram_cell[     715] = 32'hcc83462f;
    ram_cell[     716] = 32'h8a9b1759;
    ram_cell[     717] = 32'h6c7f7c40;
    ram_cell[     718] = 32'he17a6b80;
    ram_cell[     719] = 32'h10174e0c;
    ram_cell[     720] = 32'hec526b49;
    ram_cell[     721] = 32'hbec57f05;
    ram_cell[     722] = 32'h74df8109;
    ram_cell[     723] = 32'h1fc9aab8;
    ram_cell[     724] = 32'hb9b9b9a1;
    ram_cell[     725] = 32'hae93ee8e;
    ram_cell[     726] = 32'hb4bccaf8;
    ram_cell[     727] = 32'hd600b13e;
    ram_cell[     728] = 32'ha737cb5d;
    ram_cell[     729] = 32'h9f162ebb;
    ram_cell[     730] = 32'hfba0a3b7;
    ram_cell[     731] = 32'h83281f0f;
    ram_cell[     732] = 32'h9dbd1276;
    ram_cell[     733] = 32'he1860b26;
    ram_cell[     734] = 32'had806347;
    ram_cell[     735] = 32'h1bd029d3;
    ram_cell[     736] = 32'hb42b43cb;
    ram_cell[     737] = 32'h09cfb93f;
    ram_cell[     738] = 32'hf26d026f;
    ram_cell[     739] = 32'hb6ec676a;
    ram_cell[     740] = 32'hc1260e9b;
    ram_cell[     741] = 32'h5b40e977;
    ram_cell[     742] = 32'h9252d3f2;
    ram_cell[     743] = 32'h2e47ec22;
    ram_cell[     744] = 32'h7a356d85;
    ram_cell[     745] = 32'h03278eb0;
    ram_cell[     746] = 32'h0266bc88;
    ram_cell[     747] = 32'h5d7dc821;
    ram_cell[     748] = 32'h2f86cad1;
    ram_cell[     749] = 32'hfb8df94a;
    ram_cell[     750] = 32'hde7cda0e;
    ram_cell[     751] = 32'h59c8c4ab;
    ram_cell[     752] = 32'h7d7b561e;
    ram_cell[     753] = 32'h02d99dc0;
    ram_cell[     754] = 32'h27de2441;
    ram_cell[     755] = 32'h3085fe14;
    ram_cell[     756] = 32'haa02d11f;
    ram_cell[     757] = 32'h7daeb51b;
    ram_cell[     758] = 32'hd6cd9971;
    ram_cell[     759] = 32'h27ed2bfa;
    ram_cell[     760] = 32'hc64a54b2;
    ram_cell[     761] = 32'heaf94ae6;
    ram_cell[     762] = 32'h93c53690;
    ram_cell[     763] = 32'h41b438a4;
    ram_cell[     764] = 32'hfb8c3658;
    ram_cell[     765] = 32'h29117ecf;
    ram_cell[     766] = 32'h6db445be;
    ram_cell[     767] = 32'hbcf5ac05;
end

endmodule

