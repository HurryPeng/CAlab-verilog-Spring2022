`timescale 1ns / 1ps
//  功能说明
    //  ID/EX.Imm 段寄存器
// 实验要求
    // 补全模块（阶段三）

module Imm_EX(
    input wire clk, bubbleE, flushE,
    input wire [31:0] imm_in,
    output reg [31:0] imm_out
    );
    
    // TODO: Complete this module

    /* FIXME: Write your code here... */

endmodule