
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h417b06d9;
    ram_cell[       1] = 32'h0;  // 32'h7643c141;
    ram_cell[       2] = 32'h0;  // 32'h549b2a60;
    ram_cell[       3] = 32'h0;  // 32'h9202c71a;
    ram_cell[       4] = 32'h0;  // 32'hc4eb331d;
    ram_cell[       5] = 32'h0;  // 32'hcc286c75;
    ram_cell[       6] = 32'h0;  // 32'hf554d19d;
    ram_cell[       7] = 32'h0;  // 32'h95e8d2f0;
    ram_cell[       8] = 32'h0;  // 32'h44599fa0;
    ram_cell[       9] = 32'h0;  // 32'h829c91c1;
    ram_cell[      10] = 32'h0;  // 32'h3458ea1b;
    ram_cell[      11] = 32'h0;  // 32'ha19fd4a9;
    ram_cell[      12] = 32'h0;  // 32'h578c1b4f;
    ram_cell[      13] = 32'h0;  // 32'h7cfecb68;
    ram_cell[      14] = 32'h0;  // 32'haba7167a;
    ram_cell[      15] = 32'h0;  // 32'hceee0771;
    ram_cell[      16] = 32'h0;  // 32'h8bb75097;
    ram_cell[      17] = 32'h0;  // 32'h8b4ac9e1;
    ram_cell[      18] = 32'h0;  // 32'hf5afb694;
    ram_cell[      19] = 32'h0;  // 32'hfe8c2eb9;
    ram_cell[      20] = 32'h0;  // 32'hb87f6f01;
    ram_cell[      21] = 32'h0;  // 32'hcd3ddebb;
    ram_cell[      22] = 32'h0;  // 32'h19c242f3;
    ram_cell[      23] = 32'h0;  // 32'h182779c7;
    ram_cell[      24] = 32'h0;  // 32'h0a168d05;
    ram_cell[      25] = 32'h0;  // 32'h8ace0944;
    ram_cell[      26] = 32'h0;  // 32'he873ed3d;
    ram_cell[      27] = 32'h0;  // 32'h0136833d;
    ram_cell[      28] = 32'h0;  // 32'had1c0bce;
    ram_cell[      29] = 32'h0;  // 32'h65388699;
    ram_cell[      30] = 32'h0;  // 32'h954b7cb4;
    ram_cell[      31] = 32'h0;  // 32'h49ce19ea;
    ram_cell[      32] = 32'h0;  // 32'h742398d8;
    ram_cell[      33] = 32'h0;  // 32'h153db957;
    ram_cell[      34] = 32'h0;  // 32'he643ce1e;
    ram_cell[      35] = 32'h0;  // 32'hbfd3ab5b;
    ram_cell[      36] = 32'h0;  // 32'h743b6669;
    ram_cell[      37] = 32'h0;  // 32'hb553a79b;
    ram_cell[      38] = 32'h0;  // 32'h7f0d1015;
    ram_cell[      39] = 32'h0;  // 32'hd035ddad;
    ram_cell[      40] = 32'h0;  // 32'h52f681bb;
    ram_cell[      41] = 32'h0;  // 32'h270276e2;
    ram_cell[      42] = 32'h0;  // 32'hc80508c6;
    ram_cell[      43] = 32'h0;  // 32'h58d2dc82;
    ram_cell[      44] = 32'h0;  // 32'hb890b232;
    ram_cell[      45] = 32'h0;  // 32'h84ad690e;
    ram_cell[      46] = 32'h0;  // 32'h23922d34;
    ram_cell[      47] = 32'h0;  // 32'h78b21119;
    ram_cell[      48] = 32'h0;  // 32'h85eab0bc;
    ram_cell[      49] = 32'h0;  // 32'h61193978;
    ram_cell[      50] = 32'h0;  // 32'he623e21a;
    ram_cell[      51] = 32'h0;  // 32'hd29af90e;
    ram_cell[      52] = 32'h0;  // 32'h7ed28c41;
    ram_cell[      53] = 32'h0;  // 32'hd59102b8;
    ram_cell[      54] = 32'h0;  // 32'h17479949;
    ram_cell[      55] = 32'h0;  // 32'h7293a135;
    ram_cell[      56] = 32'h0;  // 32'h14ebbc91;
    ram_cell[      57] = 32'h0;  // 32'h5c09e5dd;
    ram_cell[      58] = 32'h0;  // 32'h52041350;
    ram_cell[      59] = 32'h0;  // 32'h29e322d4;
    ram_cell[      60] = 32'h0;  // 32'he4daca63;
    ram_cell[      61] = 32'h0;  // 32'hff005e7c;
    ram_cell[      62] = 32'h0;  // 32'hb2680785;
    ram_cell[      63] = 32'h0;  // 32'hd41499d4;
    ram_cell[      64] = 32'h0;  // 32'h4d44139e;
    ram_cell[      65] = 32'h0;  // 32'h3e34266e;
    ram_cell[      66] = 32'h0;  // 32'hcc650c1c;
    ram_cell[      67] = 32'h0;  // 32'h58e663c1;
    ram_cell[      68] = 32'h0;  // 32'hda1fba30;
    ram_cell[      69] = 32'h0;  // 32'he39a7016;
    ram_cell[      70] = 32'h0;  // 32'h467cfa72;
    ram_cell[      71] = 32'h0;  // 32'hffd44e23;
    ram_cell[      72] = 32'h0;  // 32'h8b75ab8b;
    ram_cell[      73] = 32'h0;  // 32'hf12e9631;
    ram_cell[      74] = 32'h0;  // 32'h70700da7;
    ram_cell[      75] = 32'h0;  // 32'h507247a1;
    ram_cell[      76] = 32'h0;  // 32'h94a745e5;
    ram_cell[      77] = 32'h0;  // 32'h62eae2fc;
    ram_cell[      78] = 32'h0;  // 32'he5f05a0d;
    ram_cell[      79] = 32'h0;  // 32'h39b3285c;
    ram_cell[      80] = 32'h0;  // 32'h2116fc4d;
    ram_cell[      81] = 32'h0;  // 32'hab5d85a6;
    ram_cell[      82] = 32'h0;  // 32'h8b84b3aa;
    ram_cell[      83] = 32'h0;  // 32'h4afda054;
    ram_cell[      84] = 32'h0;  // 32'h6f718491;
    ram_cell[      85] = 32'h0;  // 32'hb1a64819;
    ram_cell[      86] = 32'h0;  // 32'he0027f7b;
    ram_cell[      87] = 32'h0;  // 32'ha0825337;
    ram_cell[      88] = 32'h0;  // 32'hc40d3060;
    ram_cell[      89] = 32'h0;  // 32'h8ed711f7;
    ram_cell[      90] = 32'h0;  // 32'h7e6c97a8;
    ram_cell[      91] = 32'h0;  // 32'h00ebd391;
    ram_cell[      92] = 32'h0;  // 32'h16472e4c;
    ram_cell[      93] = 32'h0;  // 32'h51eb99af;
    ram_cell[      94] = 32'h0;  // 32'h103d1c0e;
    ram_cell[      95] = 32'h0;  // 32'h784427a8;
    ram_cell[      96] = 32'h0;  // 32'h6d227b09;
    ram_cell[      97] = 32'h0;  // 32'h5cd85c3d;
    ram_cell[      98] = 32'h0;  // 32'h44b09fa7;
    ram_cell[      99] = 32'h0;  // 32'hd2a2bd14;
    ram_cell[     100] = 32'h0;  // 32'h05d0bc8a;
    ram_cell[     101] = 32'h0;  // 32'h592f94da;
    ram_cell[     102] = 32'h0;  // 32'h698bb442;
    ram_cell[     103] = 32'h0;  // 32'h035cf109;
    ram_cell[     104] = 32'h0;  // 32'h2a048753;
    ram_cell[     105] = 32'h0;  // 32'hd15cda8f;
    ram_cell[     106] = 32'h0;  // 32'hb11e8fe6;
    ram_cell[     107] = 32'h0;  // 32'hcc504c5a;
    ram_cell[     108] = 32'h0;  // 32'h70935b25;
    ram_cell[     109] = 32'h0;  // 32'h2f8b82c4;
    ram_cell[     110] = 32'h0;  // 32'hfd63cf35;
    ram_cell[     111] = 32'h0;  // 32'h55b65054;
    ram_cell[     112] = 32'h0;  // 32'hc4129984;
    ram_cell[     113] = 32'h0;  // 32'haddee9de;
    ram_cell[     114] = 32'h0;  // 32'h29928731;
    ram_cell[     115] = 32'h0;  // 32'hb0192a5f;
    ram_cell[     116] = 32'h0;  // 32'h2076c5c0;
    ram_cell[     117] = 32'h0;  // 32'ha6ab229c;
    ram_cell[     118] = 32'h0;  // 32'h7eea882a;
    ram_cell[     119] = 32'h0;  // 32'ha7cb7873;
    ram_cell[     120] = 32'h0;  // 32'hd132f50e;
    ram_cell[     121] = 32'h0;  // 32'h2585af92;
    ram_cell[     122] = 32'h0;  // 32'h6ab53a90;
    ram_cell[     123] = 32'h0;  // 32'h9dc7e6c4;
    ram_cell[     124] = 32'h0;  // 32'h72692a62;
    ram_cell[     125] = 32'h0;  // 32'h3c2226d7;
    ram_cell[     126] = 32'h0;  // 32'ha63be3f3;
    ram_cell[     127] = 32'h0;  // 32'h1219357c;
    ram_cell[     128] = 32'h0;  // 32'h1ac5e72c;
    ram_cell[     129] = 32'h0;  // 32'h0ce9d676;
    ram_cell[     130] = 32'h0;  // 32'h0015d464;
    ram_cell[     131] = 32'h0;  // 32'h00347d6a;
    ram_cell[     132] = 32'h0;  // 32'h83284ea3;
    ram_cell[     133] = 32'h0;  // 32'hfd2ab52f;
    ram_cell[     134] = 32'h0;  // 32'h606d28f2;
    ram_cell[     135] = 32'h0;  // 32'h6c0850da;
    ram_cell[     136] = 32'h0;  // 32'h072559a8;
    ram_cell[     137] = 32'h0;  // 32'h6c245a9d;
    ram_cell[     138] = 32'h0;  // 32'h6295d842;
    ram_cell[     139] = 32'h0;  // 32'h10ceabbd;
    ram_cell[     140] = 32'h0;  // 32'hfeb7dfa0;
    ram_cell[     141] = 32'h0;  // 32'h55f090a5;
    ram_cell[     142] = 32'h0;  // 32'hc79e58ae;
    ram_cell[     143] = 32'h0;  // 32'hb3631345;
    ram_cell[     144] = 32'h0;  // 32'hd517b6df;
    ram_cell[     145] = 32'h0;  // 32'h24a5e5e2;
    ram_cell[     146] = 32'h0;  // 32'h3ca3a933;
    ram_cell[     147] = 32'h0;  // 32'h639dd2b3;
    ram_cell[     148] = 32'h0;  // 32'h0ed0bf8e;
    ram_cell[     149] = 32'h0;  // 32'h42f3c691;
    ram_cell[     150] = 32'h0;  // 32'h4c5829fc;
    ram_cell[     151] = 32'h0;  // 32'h99a14e2c;
    ram_cell[     152] = 32'h0;  // 32'hb72ac0ab;
    ram_cell[     153] = 32'h0;  // 32'h26d169aa;
    ram_cell[     154] = 32'h0;  // 32'hf8f6ac60;
    ram_cell[     155] = 32'h0;  // 32'h7687c6c6;
    ram_cell[     156] = 32'h0;  // 32'h6321bd0a;
    ram_cell[     157] = 32'h0;  // 32'hc5285097;
    ram_cell[     158] = 32'h0;  // 32'hd72702cd;
    ram_cell[     159] = 32'h0;  // 32'h31a53642;
    ram_cell[     160] = 32'h0;  // 32'hd05059eb;
    ram_cell[     161] = 32'h0;  // 32'hae1e12df;
    ram_cell[     162] = 32'h0;  // 32'hd4428d18;
    ram_cell[     163] = 32'h0;  // 32'hdc726681;
    ram_cell[     164] = 32'h0;  // 32'h219bf778;
    ram_cell[     165] = 32'h0;  // 32'hf12cb3c4;
    ram_cell[     166] = 32'h0;  // 32'h56dace23;
    ram_cell[     167] = 32'h0;  // 32'h062bae53;
    ram_cell[     168] = 32'h0;  // 32'h90795a63;
    ram_cell[     169] = 32'h0;  // 32'hd4a5a1b6;
    ram_cell[     170] = 32'h0;  // 32'h0cb675b2;
    ram_cell[     171] = 32'h0;  // 32'h5bb13176;
    ram_cell[     172] = 32'h0;  // 32'h18859fb6;
    ram_cell[     173] = 32'h0;  // 32'hab55e5eb;
    ram_cell[     174] = 32'h0;  // 32'h49c1fb67;
    ram_cell[     175] = 32'h0;  // 32'hd26b2128;
    ram_cell[     176] = 32'h0;  // 32'h02a51426;
    ram_cell[     177] = 32'h0;  // 32'h1c7351ac;
    ram_cell[     178] = 32'h0;  // 32'h29c085d2;
    ram_cell[     179] = 32'h0;  // 32'h54e26c52;
    ram_cell[     180] = 32'h0;  // 32'h9e5423c4;
    ram_cell[     181] = 32'h0;  // 32'h5f1c97ca;
    ram_cell[     182] = 32'h0;  // 32'h5fcf9976;
    ram_cell[     183] = 32'h0;  // 32'hc9aeea40;
    ram_cell[     184] = 32'h0;  // 32'hdc2ee53f;
    ram_cell[     185] = 32'h0;  // 32'hddf588b6;
    ram_cell[     186] = 32'h0;  // 32'haf183fc7;
    ram_cell[     187] = 32'h0;  // 32'h39877a6a;
    ram_cell[     188] = 32'h0;  // 32'hea2b9846;
    ram_cell[     189] = 32'h0;  // 32'h12189dd3;
    ram_cell[     190] = 32'h0;  // 32'h7b4c3aec;
    ram_cell[     191] = 32'h0;  // 32'h5b44e0ee;
    ram_cell[     192] = 32'h0;  // 32'hd86186bd;
    ram_cell[     193] = 32'h0;  // 32'ha0ed30b3;
    ram_cell[     194] = 32'h0;  // 32'hc02428f9;
    ram_cell[     195] = 32'h0;  // 32'hd97f7846;
    ram_cell[     196] = 32'h0;  // 32'h01c161ab;
    ram_cell[     197] = 32'h0;  // 32'ha58dd5fd;
    ram_cell[     198] = 32'h0;  // 32'h5b7ac316;
    ram_cell[     199] = 32'h0;  // 32'h1c129cf9;
    ram_cell[     200] = 32'h0;  // 32'h4f41339f;
    ram_cell[     201] = 32'h0;  // 32'h75fb943d;
    ram_cell[     202] = 32'h0;  // 32'ha9282164;
    ram_cell[     203] = 32'h0;  // 32'hc5d7c341;
    ram_cell[     204] = 32'h0;  // 32'h2398f490;
    ram_cell[     205] = 32'h0;  // 32'h2f6d37b3;
    ram_cell[     206] = 32'h0;  // 32'h56513b90;
    ram_cell[     207] = 32'h0;  // 32'hf3ca56ba;
    ram_cell[     208] = 32'h0;  // 32'he823992c;
    ram_cell[     209] = 32'h0;  // 32'hcf7155ac;
    ram_cell[     210] = 32'h0;  // 32'ha0589d69;
    ram_cell[     211] = 32'h0;  // 32'h8fe9b624;
    ram_cell[     212] = 32'h0;  // 32'hcc5ddd60;
    ram_cell[     213] = 32'h0;  // 32'ha2a96cb1;
    ram_cell[     214] = 32'h0;  // 32'h27872429;
    ram_cell[     215] = 32'h0;  // 32'h2a38f1ed;
    ram_cell[     216] = 32'h0;  // 32'hbee1efe6;
    ram_cell[     217] = 32'h0;  // 32'hb5c80b32;
    ram_cell[     218] = 32'h0;  // 32'h40990ee9;
    ram_cell[     219] = 32'h0;  // 32'h64e42d47;
    ram_cell[     220] = 32'h0;  // 32'h9eaafacf;
    ram_cell[     221] = 32'h0;  // 32'hc2e430e2;
    ram_cell[     222] = 32'h0;  // 32'hc331da46;
    ram_cell[     223] = 32'h0;  // 32'haf9d1666;
    ram_cell[     224] = 32'h0;  // 32'h870b0514;
    ram_cell[     225] = 32'h0;  // 32'h6685caf8;
    ram_cell[     226] = 32'h0;  // 32'hd4347b96;
    ram_cell[     227] = 32'h0;  // 32'h2d2e92db;
    ram_cell[     228] = 32'h0;  // 32'h08e3785c;
    ram_cell[     229] = 32'h0;  // 32'h9b81c99a;
    ram_cell[     230] = 32'h0;  // 32'hd8de19bd;
    ram_cell[     231] = 32'h0;  // 32'h7f7fa649;
    ram_cell[     232] = 32'h0;  // 32'hbd77e13a;
    ram_cell[     233] = 32'h0;  // 32'ha78241e0;
    ram_cell[     234] = 32'h0;  // 32'hd416349f;
    ram_cell[     235] = 32'h0;  // 32'hb11a1fe0;
    ram_cell[     236] = 32'h0;  // 32'h7dbcd911;
    ram_cell[     237] = 32'h0;  // 32'hb9347e65;
    ram_cell[     238] = 32'h0;  // 32'h370f7ff9;
    ram_cell[     239] = 32'h0;  // 32'h96e17637;
    ram_cell[     240] = 32'h0;  // 32'h32bf2d3c;
    ram_cell[     241] = 32'h0;  // 32'h141b5c94;
    ram_cell[     242] = 32'h0;  // 32'h6afc8311;
    ram_cell[     243] = 32'h0;  // 32'h953f32f1;
    ram_cell[     244] = 32'h0;  // 32'ha168383e;
    ram_cell[     245] = 32'h0;  // 32'h83e9804a;
    ram_cell[     246] = 32'h0;  // 32'h0e60beab;
    ram_cell[     247] = 32'h0;  // 32'h46d924c1;
    ram_cell[     248] = 32'h0;  // 32'h21b39c36;
    ram_cell[     249] = 32'h0;  // 32'h7551df1f;
    ram_cell[     250] = 32'h0;  // 32'hf0c2763a;
    ram_cell[     251] = 32'h0;  // 32'h1d0f26c1;
    ram_cell[     252] = 32'h0;  // 32'h024ad7d3;
    ram_cell[     253] = 32'h0;  // 32'h400f973a;
    ram_cell[     254] = 32'h0;  // 32'hfd5d63ce;
    ram_cell[     255] = 32'h0;  // 32'hd0e7e463;
    // src matrix A
    ram_cell[     256] = 32'hb8ae64d2;
    ram_cell[     257] = 32'h5b85b124;
    ram_cell[     258] = 32'hf1a99349;
    ram_cell[     259] = 32'h7a6de1d3;
    ram_cell[     260] = 32'hd96d7019;
    ram_cell[     261] = 32'he6f5c05c;
    ram_cell[     262] = 32'h765f2fc3;
    ram_cell[     263] = 32'hee7b742d;
    ram_cell[     264] = 32'h858fbc38;
    ram_cell[     265] = 32'he2e54dcc;
    ram_cell[     266] = 32'ha7c812c0;
    ram_cell[     267] = 32'h50508da9;
    ram_cell[     268] = 32'h47ad541a;
    ram_cell[     269] = 32'h400828f7;
    ram_cell[     270] = 32'h19fb5c31;
    ram_cell[     271] = 32'h9ae98948;
    ram_cell[     272] = 32'ha4e0522a;
    ram_cell[     273] = 32'hc1e1a79f;
    ram_cell[     274] = 32'haf686ac6;
    ram_cell[     275] = 32'h0c699d91;
    ram_cell[     276] = 32'h6aae34b8;
    ram_cell[     277] = 32'hadf71ef5;
    ram_cell[     278] = 32'h9a9c9b01;
    ram_cell[     279] = 32'hbd9788f4;
    ram_cell[     280] = 32'hfa3e6d96;
    ram_cell[     281] = 32'hba08508c;
    ram_cell[     282] = 32'h4688a20d;
    ram_cell[     283] = 32'he36b5b0c;
    ram_cell[     284] = 32'h341dceb7;
    ram_cell[     285] = 32'h3a766b58;
    ram_cell[     286] = 32'he045f235;
    ram_cell[     287] = 32'he1164f16;
    ram_cell[     288] = 32'hd3824311;
    ram_cell[     289] = 32'h6b817c93;
    ram_cell[     290] = 32'hf22e460c;
    ram_cell[     291] = 32'h1776a0d4;
    ram_cell[     292] = 32'h6796ef62;
    ram_cell[     293] = 32'h7704bb57;
    ram_cell[     294] = 32'h5aaffaeb;
    ram_cell[     295] = 32'h7e7d02b1;
    ram_cell[     296] = 32'haf7fc57f;
    ram_cell[     297] = 32'h89e1c9e0;
    ram_cell[     298] = 32'h3bdd782b;
    ram_cell[     299] = 32'h7ca4b688;
    ram_cell[     300] = 32'h745d4685;
    ram_cell[     301] = 32'hb26dc44a;
    ram_cell[     302] = 32'hc5d1dd2c;
    ram_cell[     303] = 32'he38442a2;
    ram_cell[     304] = 32'h9e1bee2f;
    ram_cell[     305] = 32'h44fc7a65;
    ram_cell[     306] = 32'h5f3a64f5;
    ram_cell[     307] = 32'h4de11ebd;
    ram_cell[     308] = 32'hfd650c1b;
    ram_cell[     309] = 32'heece378a;
    ram_cell[     310] = 32'h22f3debf;
    ram_cell[     311] = 32'he3f67a28;
    ram_cell[     312] = 32'hfe221688;
    ram_cell[     313] = 32'he829c05f;
    ram_cell[     314] = 32'hc40edd72;
    ram_cell[     315] = 32'h9ea5a406;
    ram_cell[     316] = 32'hb079cada;
    ram_cell[     317] = 32'h50ee2d02;
    ram_cell[     318] = 32'hc6f7add3;
    ram_cell[     319] = 32'hc9c119fa;
    ram_cell[     320] = 32'h4115b59e;
    ram_cell[     321] = 32'hcaea928d;
    ram_cell[     322] = 32'h7681ea3f;
    ram_cell[     323] = 32'h89ba5bb3;
    ram_cell[     324] = 32'hea66a493;
    ram_cell[     325] = 32'he67a8239;
    ram_cell[     326] = 32'he87ad50b;
    ram_cell[     327] = 32'hfd19b9ab;
    ram_cell[     328] = 32'hb2318817;
    ram_cell[     329] = 32'h32d2e0ee;
    ram_cell[     330] = 32'hccadac4e;
    ram_cell[     331] = 32'h47667293;
    ram_cell[     332] = 32'h89967dc0;
    ram_cell[     333] = 32'h586f21a7;
    ram_cell[     334] = 32'h98b64d8c;
    ram_cell[     335] = 32'h8c42fe5c;
    ram_cell[     336] = 32'he018479b;
    ram_cell[     337] = 32'h4ab20883;
    ram_cell[     338] = 32'hc8defd1f;
    ram_cell[     339] = 32'hb092a905;
    ram_cell[     340] = 32'hd5687d56;
    ram_cell[     341] = 32'hb84b693e;
    ram_cell[     342] = 32'h351722ce;
    ram_cell[     343] = 32'h6fff1024;
    ram_cell[     344] = 32'h6ed3c675;
    ram_cell[     345] = 32'hfc82e514;
    ram_cell[     346] = 32'hf66b8662;
    ram_cell[     347] = 32'hac2ae151;
    ram_cell[     348] = 32'h101f6dfe;
    ram_cell[     349] = 32'h46906b7f;
    ram_cell[     350] = 32'hce99f7c7;
    ram_cell[     351] = 32'hd0dbb4cd;
    ram_cell[     352] = 32'hc3db3571;
    ram_cell[     353] = 32'ha0c442b5;
    ram_cell[     354] = 32'h2a7be809;
    ram_cell[     355] = 32'h0956103d;
    ram_cell[     356] = 32'hfca82c33;
    ram_cell[     357] = 32'h4cb6c7d4;
    ram_cell[     358] = 32'he413c086;
    ram_cell[     359] = 32'hccd42479;
    ram_cell[     360] = 32'h3c429b25;
    ram_cell[     361] = 32'hed279201;
    ram_cell[     362] = 32'hfef4d0f4;
    ram_cell[     363] = 32'he8152a43;
    ram_cell[     364] = 32'h885a35f1;
    ram_cell[     365] = 32'hbb962447;
    ram_cell[     366] = 32'hf1fc1371;
    ram_cell[     367] = 32'hc1259015;
    ram_cell[     368] = 32'h6c6c0bcf;
    ram_cell[     369] = 32'ha0628c70;
    ram_cell[     370] = 32'h60892a12;
    ram_cell[     371] = 32'h5ed14659;
    ram_cell[     372] = 32'hcef30263;
    ram_cell[     373] = 32'h1c52c780;
    ram_cell[     374] = 32'h4e23b2d1;
    ram_cell[     375] = 32'h0a6a1d5d;
    ram_cell[     376] = 32'h421833a6;
    ram_cell[     377] = 32'h44ba0a5b;
    ram_cell[     378] = 32'h65780874;
    ram_cell[     379] = 32'h370274c5;
    ram_cell[     380] = 32'h9fe15828;
    ram_cell[     381] = 32'h469db72e;
    ram_cell[     382] = 32'hb4cd2e85;
    ram_cell[     383] = 32'hb29f5d04;
    ram_cell[     384] = 32'h85bebdc6;
    ram_cell[     385] = 32'h34671c7f;
    ram_cell[     386] = 32'h5b013648;
    ram_cell[     387] = 32'h3eeb52f0;
    ram_cell[     388] = 32'h5793726c;
    ram_cell[     389] = 32'h5651fbb8;
    ram_cell[     390] = 32'h9792288d;
    ram_cell[     391] = 32'h784e2740;
    ram_cell[     392] = 32'h2e48c5fb;
    ram_cell[     393] = 32'h4a8a3938;
    ram_cell[     394] = 32'h680b24fd;
    ram_cell[     395] = 32'hfa5ad918;
    ram_cell[     396] = 32'h242bfcd5;
    ram_cell[     397] = 32'h810a48f0;
    ram_cell[     398] = 32'h5657eadb;
    ram_cell[     399] = 32'he70ee4cd;
    ram_cell[     400] = 32'hb3259352;
    ram_cell[     401] = 32'heb7b27e8;
    ram_cell[     402] = 32'h9e5d1f2d;
    ram_cell[     403] = 32'h96b2adb3;
    ram_cell[     404] = 32'h5efd9752;
    ram_cell[     405] = 32'h38c11e52;
    ram_cell[     406] = 32'h86fcd9a6;
    ram_cell[     407] = 32'h31d18a9c;
    ram_cell[     408] = 32'h7bd5d2e0;
    ram_cell[     409] = 32'he5920ecf;
    ram_cell[     410] = 32'hd9bef594;
    ram_cell[     411] = 32'h1d83b5ba;
    ram_cell[     412] = 32'h67bf278d;
    ram_cell[     413] = 32'h4f9435c2;
    ram_cell[     414] = 32'h1a433d02;
    ram_cell[     415] = 32'h89a7a8c0;
    ram_cell[     416] = 32'h74b81df9;
    ram_cell[     417] = 32'h6ecd90f5;
    ram_cell[     418] = 32'h1f82ee79;
    ram_cell[     419] = 32'h2e5f0d98;
    ram_cell[     420] = 32'h9ef3ee5c;
    ram_cell[     421] = 32'hd1626887;
    ram_cell[     422] = 32'h1da482df;
    ram_cell[     423] = 32'h058d9825;
    ram_cell[     424] = 32'hff79824f;
    ram_cell[     425] = 32'h09813ef7;
    ram_cell[     426] = 32'h47b168ba;
    ram_cell[     427] = 32'he1d1fb1c;
    ram_cell[     428] = 32'hfae129f2;
    ram_cell[     429] = 32'h76eb67db;
    ram_cell[     430] = 32'hb75dfdf8;
    ram_cell[     431] = 32'h9035cd9c;
    ram_cell[     432] = 32'he7180b4f;
    ram_cell[     433] = 32'hafa5846e;
    ram_cell[     434] = 32'h5c7cbe45;
    ram_cell[     435] = 32'hb057be5e;
    ram_cell[     436] = 32'h64df4394;
    ram_cell[     437] = 32'h9b2be037;
    ram_cell[     438] = 32'hf6569969;
    ram_cell[     439] = 32'he4582ea6;
    ram_cell[     440] = 32'hc73890bf;
    ram_cell[     441] = 32'h37fe6f7b;
    ram_cell[     442] = 32'ha57960b3;
    ram_cell[     443] = 32'hafae0b72;
    ram_cell[     444] = 32'h8bd4b8e4;
    ram_cell[     445] = 32'h8346df6b;
    ram_cell[     446] = 32'hfc800ff9;
    ram_cell[     447] = 32'hf0ae7730;
    ram_cell[     448] = 32'he4e2a3a5;
    ram_cell[     449] = 32'h8054f706;
    ram_cell[     450] = 32'h82f9af5e;
    ram_cell[     451] = 32'hfa1ef5e6;
    ram_cell[     452] = 32'h8176bee7;
    ram_cell[     453] = 32'hf94aa04f;
    ram_cell[     454] = 32'hbb4459ab;
    ram_cell[     455] = 32'h90df3027;
    ram_cell[     456] = 32'h81ff5707;
    ram_cell[     457] = 32'h58cc6211;
    ram_cell[     458] = 32'h13f408a4;
    ram_cell[     459] = 32'hd7370140;
    ram_cell[     460] = 32'h898651dc;
    ram_cell[     461] = 32'h3eb31ea7;
    ram_cell[     462] = 32'h95da4af0;
    ram_cell[     463] = 32'hb5c283f7;
    ram_cell[     464] = 32'h7f3b3b20;
    ram_cell[     465] = 32'h758b2e4c;
    ram_cell[     466] = 32'he9aa0acf;
    ram_cell[     467] = 32'h6190b632;
    ram_cell[     468] = 32'h0164bcbb;
    ram_cell[     469] = 32'h06a1412d;
    ram_cell[     470] = 32'h44c803e1;
    ram_cell[     471] = 32'hd3b96234;
    ram_cell[     472] = 32'hd963c5c1;
    ram_cell[     473] = 32'hc7517b04;
    ram_cell[     474] = 32'he76bde6d;
    ram_cell[     475] = 32'h453d3730;
    ram_cell[     476] = 32'h5b4a4e4a;
    ram_cell[     477] = 32'h4b9c8edb;
    ram_cell[     478] = 32'hdda335dc;
    ram_cell[     479] = 32'h67515079;
    ram_cell[     480] = 32'hd4fb4f7a;
    ram_cell[     481] = 32'h93231156;
    ram_cell[     482] = 32'he2dfd007;
    ram_cell[     483] = 32'h54b446c4;
    ram_cell[     484] = 32'h34c661b9;
    ram_cell[     485] = 32'hd03b9918;
    ram_cell[     486] = 32'hc03df8ac;
    ram_cell[     487] = 32'h1707b1df;
    ram_cell[     488] = 32'h91c7c56f;
    ram_cell[     489] = 32'hb96b33d6;
    ram_cell[     490] = 32'hd39a7110;
    ram_cell[     491] = 32'h0390e88a;
    ram_cell[     492] = 32'h8698719d;
    ram_cell[     493] = 32'h95b5fe2a;
    ram_cell[     494] = 32'h3763f9a0;
    ram_cell[     495] = 32'h7b4cf7d5;
    ram_cell[     496] = 32'h2874cf5a;
    ram_cell[     497] = 32'he004c5e0;
    ram_cell[     498] = 32'h637b6b53;
    ram_cell[     499] = 32'h119ebc92;
    ram_cell[     500] = 32'h87794ee1;
    ram_cell[     501] = 32'h6ef4a58f;
    ram_cell[     502] = 32'hf353d326;
    ram_cell[     503] = 32'ha2861a40;
    ram_cell[     504] = 32'he87cc643;
    ram_cell[     505] = 32'h441526ec;
    ram_cell[     506] = 32'hfaae948f;
    ram_cell[     507] = 32'h774f92d7;
    ram_cell[     508] = 32'h35fc1718;
    ram_cell[     509] = 32'hb7adcebe;
    ram_cell[     510] = 32'h3062fb99;
    ram_cell[     511] = 32'h96a48aa9;
    // src matrix B
    ram_cell[     512] = 32'h27ccb18f;
    ram_cell[     513] = 32'h393900c4;
    ram_cell[     514] = 32'h54855a13;
    ram_cell[     515] = 32'h4c988ac1;
    ram_cell[     516] = 32'he27422f1;
    ram_cell[     517] = 32'hef88ea0f;
    ram_cell[     518] = 32'hccd2e53e;
    ram_cell[     519] = 32'h2601f5be;
    ram_cell[     520] = 32'hd667e07a;
    ram_cell[     521] = 32'h16d1d61b;
    ram_cell[     522] = 32'hee495498;
    ram_cell[     523] = 32'hd4ee6bd5;
    ram_cell[     524] = 32'h0a2e0b07;
    ram_cell[     525] = 32'h3ef1812d;
    ram_cell[     526] = 32'h01a6e7da;
    ram_cell[     527] = 32'h8ade6f50;
    ram_cell[     528] = 32'h4aad786d;
    ram_cell[     529] = 32'h45cc6f60;
    ram_cell[     530] = 32'h457e18d5;
    ram_cell[     531] = 32'hd0447f44;
    ram_cell[     532] = 32'h3643c3e7;
    ram_cell[     533] = 32'hb4e1e915;
    ram_cell[     534] = 32'h02ca2d22;
    ram_cell[     535] = 32'he292112c;
    ram_cell[     536] = 32'h8f7b97e4;
    ram_cell[     537] = 32'h1a77b578;
    ram_cell[     538] = 32'h38dfed0b;
    ram_cell[     539] = 32'h4e6682a3;
    ram_cell[     540] = 32'hb3af922a;
    ram_cell[     541] = 32'h9243ad6f;
    ram_cell[     542] = 32'ha1824997;
    ram_cell[     543] = 32'hb89bf489;
    ram_cell[     544] = 32'he3480148;
    ram_cell[     545] = 32'h08f4cfb2;
    ram_cell[     546] = 32'h4c218d90;
    ram_cell[     547] = 32'hc50d5652;
    ram_cell[     548] = 32'hc76c3aac;
    ram_cell[     549] = 32'h43187a50;
    ram_cell[     550] = 32'h8109fcdc;
    ram_cell[     551] = 32'hfa8f39a1;
    ram_cell[     552] = 32'h29c464f6;
    ram_cell[     553] = 32'h9f3d0d76;
    ram_cell[     554] = 32'hbefc74af;
    ram_cell[     555] = 32'h5db62b72;
    ram_cell[     556] = 32'h579463f0;
    ram_cell[     557] = 32'h72dc9292;
    ram_cell[     558] = 32'he6dd1445;
    ram_cell[     559] = 32'h29187ad2;
    ram_cell[     560] = 32'h3843baf3;
    ram_cell[     561] = 32'hfeabc225;
    ram_cell[     562] = 32'h0b12518a;
    ram_cell[     563] = 32'hd3a062f5;
    ram_cell[     564] = 32'hb5703edf;
    ram_cell[     565] = 32'h7c934243;
    ram_cell[     566] = 32'he237b46d;
    ram_cell[     567] = 32'h1852f0ed;
    ram_cell[     568] = 32'hfcf539c6;
    ram_cell[     569] = 32'h11b9185d;
    ram_cell[     570] = 32'h254ea1cd;
    ram_cell[     571] = 32'hef37b9bb;
    ram_cell[     572] = 32'hd3a8a10f;
    ram_cell[     573] = 32'h0c237b31;
    ram_cell[     574] = 32'hc6b90713;
    ram_cell[     575] = 32'hc01611da;
    ram_cell[     576] = 32'h68d80da1;
    ram_cell[     577] = 32'hbe069c81;
    ram_cell[     578] = 32'h543b5ae4;
    ram_cell[     579] = 32'h374c6467;
    ram_cell[     580] = 32'hb6901904;
    ram_cell[     581] = 32'h50c4262b;
    ram_cell[     582] = 32'h0b163af5;
    ram_cell[     583] = 32'h4df64668;
    ram_cell[     584] = 32'h3821ac9e;
    ram_cell[     585] = 32'hcd5a1a24;
    ram_cell[     586] = 32'h6be1a39d;
    ram_cell[     587] = 32'hf46970f2;
    ram_cell[     588] = 32'he0b4dda9;
    ram_cell[     589] = 32'ha72327f0;
    ram_cell[     590] = 32'h8601e442;
    ram_cell[     591] = 32'h7b58ad4c;
    ram_cell[     592] = 32'h96f72384;
    ram_cell[     593] = 32'h5f4d9cb3;
    ram_cell[     594] = 32'hfc557c64;
    ram_cell[     595] = 32'h414d627c;
    ram_cell[     596] = 32'h2c79b28a;
    ram_cell[     597] = 32'he77454a4;
    ram_cell[     598] = 32'h10e0ba79;
    ram_cell[     599] = 32'h1cd6b298;
    ram_cell[     600] = 32'h0885a3cd;
    ram_cell[     601] = 32'hfdfd48a5;
    ram_cell[     602] = 32'h494df440;
    ram_cell[     603] = 32'ha530d65e;
    ram_cell[     604] = 32'hd2c99b45;
    ram_cell[     605] = 32'h6fbec9e1;
    ram_cell[     606] = 32'h2e93de7b;
    ram_cell[     607] = 32'h9a77bd99;
    ram_cell[     608] = 32'h404df4ea;
    ram_cell[     609] = 32'h2fa364f2;
    ram_cell[     610] = 32'h9f91b19c;
    ram_cell[     611] = 32'hbd05babd;
    ram_cell[     612] = 32'h20a69ab9;
    ram_cell[     613] = 32'h3d16e750;
    ram_cell[     614] = 32'hf42a8283;
    ram_cell[     615] = 32'h8a8165eb;
    ram_cell[     616] = 32'hce6e24fc;
    ram_cell[     617] = 32'h3c6c388f;
    ram_cell[     618] = 32'hcf991908;
    ram_cell[     619] = 32'h51a0b87b;
    ram_cell[     620] = 32'h04d445b8;
    ram_cell[     621] = 32'hc71a7548;
    ram_cell[     622] = 32'he333c583;
    ram_cell[     623] = 32'hf31e6828;
    ram_cell[     624] = 32'ha73cfc89;
    ram_cell[     625] = 32'hce7d8eaf;
    ram_cell[     626] = 32'h761b0b6e;
    ram_cell[     627] = 32'hd0682767;
    ram_cell[     628] = 32'h6338aebc;
    ram_cell[     629] = 32'h81b4ed26;
    ram_cell[     630] = 32'h4d677d17;
    ram_cell[     631] = 32'hb772bdc2;
    ram_cell[     632] = 32'h3c69fa84;
    ram_cell[     633] = 32'ha3f744ab;
    ram_cell[     634] = 32'he64f7701;
    ram_cell[     635] = 32'h865e8260;
    ram_cell[     636] = 32'h382f6069;
    ram_cell[     637] = 32'hbcfeed33;
    ram_cell[     638] = 32'hf2209f04;
    ram_cell[     639] = 32'h9f21c238;
    ram_cell[     640] = 32'h3d0d4dea;
    ram_cell[     641] = 32'h75b4fae0;
    ram_cell[     642] = 32'hd873add8;
    ram_cell[     643] = 32'hbf62b1c4;
    ram_cell[     644] = 32'he3bd1d8b;
    ram_cell[     645] = 32'hd5345b96;
    ram_cell[     646] = 32'h663c4773;
    ram_cell[     647] = 32'h64f36ec5;
    ram_cell[     648] = 32'h89090aee;
    ram_cell[     649] = 32'h16325234;
    ram_cell[     650] = 32'h0fb885d1;
    ram_cell[     651] = 32'hb3fff2c1;
    ram_cell[     652] = 32'h5347c5a9;
    ram_cell[     653] = 32'he19567d1;
    ram_cell[     654] = 32'hf1c86eb1;
    ram_cell[     655] = 32'h63074ef7;
    ram_cell[     656] = 32'hfc7214c4;
    ram_cell[     657] = 32'h21207a6c;
    ram_cell[     658] = 32'h57c806c1;
    ram_cell[     659] = 32'h21847e77;
    ram_cell[     660] = 32'hc20be3ae;
    ram_cell[     661] = 32'h0644a7bc;
    ram_cell[     662] = 32'h485235ed;
    ram_cell[     663] = 32'hf497b38c;
    ram_cell[     664] = 32'hde2ff963;
    ram_cell[     665] = 32'hd86cd8c3;
    ram_cell[     666] = 32'h16eede10;
    ram_cell[     667] = 32'h5ce9ca7e;
    ram_cell[     668] = 32'hb1eb7c36;
    ram_cell[     669] = 32'h1614c00c;
    ram_cell[     670] = 32'h1ca5187d;
    ram_cell[     671] = 32'hee25136f;
    ram_cell[     672] = 32'h404d1049;
    ram_cell[     673] = 32'h344488fe;
    ram_cell[     674] = 32'hab83d282;
    ram_cell[     675] = 32'h7b9c497b;
    ram_cell[     676] = 32'h0aaa11aa;
    ram_cell[     677] = 32'h5f272a43;
    ram_cell[     678] = 32'h503d10bb;
    ram_cell[     679] = 32'h65acb4e7;
    ram_cell[     680] = 32'hff99f53a;
    ram_cell[     681] = 32'hdcce8ac4;
    ram_cell[     682] = 32'haf2ba485;
    ram_cell[     683] = 32'hef90b83b;
    ram_cell[     684] = 32'hf7976fe1;
    ram_cell[     685] = 32'hd9e7c84b;
    ram_cell[     686] = 32'h3ffa5b30;
    ram_cell[     687] = 32'h77bc2ab7;
    ram_cell[     688] = 32'hc9c1bf2e;
    ram_cell[     689] = 32'h6ec35ec1;
    ram_cell[     690] = 32'hfd71c9ce;
    ram_cell[     691] = 32'h28a41fe4;
    ram_cell[     692] = 32'h8acb8b54;
    ram_cell[     693] = 32'hc74e2771;
    ram_cell[     694] = 32'h5761ab6e;
    ram_cell[     695] = 32'hb10dcda9;
    ram_cell[     696] = 32'h4a44421d;
    ram_cell[     697] = 32'h0cc95b38;
    ram_cell[     698] = 32'hd2d59c81;
    ram_cell[     699] = 32'hdada6e93;
    ram_cell[     700] = 32'h2ea79164;
    ram_cell[     701] = 32'ha69460d1;
    ram_cell[     702] = 32'h7710e982;
    ram_cell[     703] = 32'ha288d5cf;
    ram_cell[     704] = 32'haeafabe0;
    ram_cell[     705] = 32'hc2589383;
    ram_cell[     706] = 32'h09471f46;
    ram_cell[     707] = 32'h849f337f;
    ram_cell[     708] = 32'h593ffcb1;
    ram_cell[     709] = 32'h677e9058;
    ram_cell[     710] = 32'h9db27fe0;
    ram_cell[     711] = 32'h27ed6286;
    ram_cell[     712] = 32'ha78cc68c;
    ram_cell[     713] = 32'ha4a35aee;
    ram_cell[     714] = 32'h5126fb84;
    ram_cell[     715] = 32'hfcef2fe9;
    ram_cell[     716] = 32'h7565f9bf;
    ram_cell[     717] = 32'h9e36b100;
    ram_cell[     718] = 32'hce7bc7d8;
    ram_cell[     719] = 32'hc274ba13;
    ram_cell[     720] = 32'hf2f2429c;
    ram_cell[     721] = 32'hd4172a69;
    ram_cell[     722] = 32'hd256a8d5;
    ram_cell[     723] = 32'h8c22020b;
    ram_cell[     724] = 32'he70a1f04;
    ram_cell[     725] = 32'hdccaf01e;
    ram_cell[     726] = 32'ha91530ec;
    ram_cell[     727] = 32'h12622b76;
    ram_cell[     728] = 32'h6d95a18f;
    ram_cell[     729] = 32'hd2d8f32b;
    ram_cell[     730] = 32'h1c560c36;
    ram_cell[     731] = 32'h6461d71a;
    ram_cell[     732] = 32'hcb241066;
    ram_cell[     733] = 32'h7a7ad944;
    ram_cell[     734] = 32'h53ef831d;
    ram_cell[     735] = 32'hacad6ac8;
    ram_cell[     736] = 32'hebf6ecae;
    ram_cell[     737] = 32'hd856d758;
    ram_cell[     738] = 32'h0e2f5c69;
    ram_cell[     739] = 32'h3256388b;
    ram_cell[     740] = 32'haae5e777;
    ram_cell[     741] = 32'he359f010;
    ram_cell[     742] = 32'h4873f7e1;
    ram_cell[     743] = 32'hb197b668;
    ram_cell[     744] = 32'ha0aa3384;
    ram_cell[     745] = 32'h74ccab8d;
    ram_cell[     746] = 32'h1be1e2e0;
    ram_cell[     747] = 32'ha0fb7536;
    ram_cell[     748] = 32'h4f7bafec;
    ram_cell[     749] = 32'h251ecae7;
    ram_cell[     750] = 32'h550952ce;
    ram_cell[     751] = 32'h150b2336;
    ram_cell[     752] = 32'hd0daf2d4;
    ram_cell[     753] = 32'h8e9c0dd7;
    ram_cell[     754] = 32'h0c91a4a2;
    ram_cell[     755] = 32'h066041b4;
    ram_cell[     756] = 32'h7a326a70;
    ram_cell[     757] = 32'h3912ae51;
    ram_cell[     758] = 32'h1b3eda58;
    ram_cell[     759] = 32'h203779ad;
    ram_cell[     760] = 32'h51c7e726;
    ram_cell[     761] = 32'hd7fe23db;
    ram_cell[     762] = 32'hf7160623;
    ram_cell[     763] = 32'hc54def20;
    ram_cell[     764] = 32'h31d540f9;
    ram_cell[     765] = 32'hd2af3ee5;
    ram_cell[     766] = 32'h4acc35e9;
    ram_cell[     767] = 32'hf7ff3865;
end

endmodule

